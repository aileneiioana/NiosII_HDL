
module HelloNiosIntr (
	clk_clk);	

	input		clk_clk;
endmodule
