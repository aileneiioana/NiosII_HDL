// nios_custom_dma.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module nios_custom_dma (
		input  wire  clk_clk  // clk.clk
	);

	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [18:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] simple_dma_read_master_readdata;                             // mm_interconnect_0:simple_dma_read_master_readdata -> simple_dma:avm_read_master_readdata
	wire         simple_dma_read_master_waitrequest;                          // mm_interconnect_0:simple_dma_read_master_waitrequest -> simple_dma:avm_read_master_waitrequest
	wire         simple_dma_read_master_read;                                 // simple_dma:avm_read_master_read -> mm_interconnect_0:simple_dma_read_master_read
	wire  [31:0] simple_dma_read_master_address;                              // simple_dma:avm_read_master_address -> mm_interconnect_0:simple_dma_read_master_address
	wire  [31:0] pipelined_dma_read_master_readdata;                          // mm_interconnect_0:pipelined_dma_read_master_readdata -> pipelined_dma:avm_read_master_readdata
	wire         pipelined_dma_read_master_waitrequest;                       // mm_interconnect_0:pipelined_dma_read_master_waitrequest -> pipelined_dma:avm_read_master_waitrequest
	wire         pipelined_dma_read_master_read;                              // pipelined_dma:avm_read_master_read -> mm_interconnect_0:pipelined_dma_read_master_read
	wire  [31:0] pipelined_dma_read_master_address;                           // pipelined_dma:avm_read_master_address -> mm_interconnect_0:pipelined_dma_read_master_address
	wire         pipelined_dma_read_master_readdatavalid;                     // mm_interconnect_0:pipelined_dma_read_master_readdatavalid -> pipelined_dma:avm_read_master_readdatavalid
	wire  [31:0] burst_dma_read_master_readdata;                              // mm_interconnect_0:burst_dma_read_master_readdata -> burst_dma:avm_read_master_readdata
	wire         burst_dma_read_master_waitrequest;                           // mm_interconnect_0:burst_dma_read_master_waitrequest -> burst_dma:avm_read_master_waitrequest
	wire         burst_dma_read_master_read;                                  // burst_dma:avm_read_master_read -> mm_interconnect_0:burst_dma_read_master_read
	wire  [31:0] burst_dma_read_master_address;                               // burst_dma:avm_read_master_address -> mm_interconnect_0:burst_dma_read_master_address
	wire         burst_dma_read_master_readdatavalid;                         // mm_interconnect_0:burst_dma_read_master_readdatavalid -> burst_dma:avm_read_master_readdatavalid
	wire   [5:0] burst_dma_read_master_burstcount;                            // burst_dma:avm_read_master_burstcount -> mm_interconnect_0:burst_dma_read_master_burstcount
	wire  [31:0] block_dma_read_master_readdata;                              // mm_interconnect_0:block_dma_read_master_readdata -> block_dma:avm_read_master_readdata
	wire         block_dma_read_master_waitrequest;                           // mm_interconnect_0:block_dma_read_master_waitrequest -> block_dma:avm_read_master_waitrequest
	wire         block_dma_read_master_read;                                  // block_dma:avm_read_master_read -> mm_interconnect_0:block_dma_read_master_read
	wire  [31:0] block_dma_read_master_address;                               // block_dma:avm_read_master_address -> mm_interconnect_0:block_dma_read_master_address
	wire         simple_dma_write_master_waitrequest;                         // mm_interconnect_0:simple_dma_write_master_waitrequest -> simple_dma:avm_write_master_waitrequest
	wire  [31:0] simple_dma_write_master_address;                             // simple_dma:avm_write_master_address -> mm_interconnect_0:simple_dma_write_master_address
	wire         simple_dma_write_master_write;                               // simple_dma:avm_write_master_write -> mm_interconnect_0:simple_dma_write_master_write
	wire  [31:0] simple_dma_write_master_writedata;                           // simple_dma:avm_write_master_writedata -> mm_interconnect_0:simple_dma_write_master_writedata
	wire         pipelined_dma_write_master_waitrequest;                      // mm_interconnect_0:pipelined_dma_write_master_waitrequest -> pipelined_dma:avm_write_master_waitrequest
	wire  [31:0] pipelined_dma_write_master_address;                          // pipelined_dma:avm_write_master_address -> mm_interconnect_0:pipelined_dma_write_master_address
	wire         pipelined_dma_write_master_write;                            // pipelined_dma:avm_write_master_write -> mm_interconnect_0:pipelined_dma_write_master_write
	wire  [31:0] pipelined_dma_write_master_writedata;                        // pipelined_dma:avm_write_master_writedata -> mm_interconnect_0:pipelined_dma_write_master_writedata
	wire         burst_dma_write_master_waitrequest;                          // mm_interconnect_0:burst_dma_write_master_waitrequest -> burst_dma:avm_write_master_waitrequest
	wire  [31:0] burst_dma_write_master_address;                              // burst_dma:avm_write_master_address -> mm_interconnect_0:burst_dma_write_master_address
	wire         burst_dma_write_master_write;                                // burst_dma:avm_write_master_write -> mm_interconnect_0:burst_dma_write_master_write
	wire  [31:0] burst_dma_write_master_writedata;                            // burst_dma:avm_write_master_writedata -> mm_interconnect_0:burst_dma_write_master_writedata
	wire   [5:0] burst_dma_write_master_burstcount;                           // burst_dma:avm_write_master_burstcount -> mm_interconnect_0:burst_dma_write_master_burstcount
	wire         block_dma_write_master_waitrequest;                          // mm_interconnect_0:block_dma_write_master_waitrequest -> block_dma:avm_write_master_waitrequest
	wire  [31:0] block_dma_write_master_address;                              // block_dma:avm_write_master_address -> mm_interconnect_0:block_dma_write_master_address
	wire         block_dma_write_master_write;                                // block_dma:avm_write_master_write -> mm_interconnect_0:block_dma_write_master_write
	wire  [31:0] block_dma_write_master_writedata;                            // block_dma:avm_write_master_writedata -> mm_interconnect_0:block_dma_write_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [18:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_simple_dma_csr_readdata;                   // simple_dma:avs_csr_readdata -> mm_interconnect_0:simple_dma_csr_readdata
	wire   [1:0] mm_interconnect_0_simple_dma_csr_address;                    // mm_interconnect_0:simple_dma_csr_address -> simple_dma:avs_csr_address
	wire         mm_interconnect_0_simple_dma_csr_write;                      // mm_interconnect_0:simple_dma_csr_write -> simple_dma:avs_csr_write
	wire  [31:0] mm_interconnect_0_simple_dma_csr_writedata;                  // mm_interconnect_0:simple_dma_csr_writedata -> simple_dma:avs_csr_writedata
	wire  [31:0] mm_interconnect_0_pipelined_dma_csr_readdata;                // pipelined_dma:avs_csr_readdata -> mm_interconnect_0:pipelined_dma_csr_readdata
	wire   [1:0] mm_interconnect_0_pipelined_dma_csr_address;                 // mm_interconnect_0:pipelined_dma_csr_address -> pipelined_dma:avs_csr_address
	wire         mm_interconnect_0_pipelined_dma_csr_write;                   // mm_interconnect_0:pipelined_dma_csr_write -> pipelined_dma:avs_csr_write
	wire  [31:0] mm_interconnect_0_pipelined_dma_csr_writedata;               // mm_interconnect_0:pipelined_dma_csr_writedata -> pipelined_dma:avs_csr_writedata
	wire  [31:0] mm_interconnect_0_burst_dma_csr_readdata;                    // burst_dma:avs_csr_readdata -> mm_interconnect_0:burst_dma_csr_readdata
	wire   [1:0] mm_interconnect_0_burst_dma_csr_address;                     // mm_interconnect_0:burst_dma_csr_address -> burst_dma:avs_csr_address
	wire         mm_interconnect_0_burst_dma_csr_write;                       // mm_interconnect_0:burst_dma_csr_write -> burst_dma:avs_csr_write
	wire  [31:0] mm_interconnect_0_burst_dma_csr_writedata;                   // mm_interconnect_0:burst_dma_csr_writedata -> burst_dma:avs_csr_writedata
	wire  [31:0] mm_interconnect_0_block_dma_csr_readdata;                    // block_dma:avs_csr_readdata -> mm_interconnect_0:block_dma_csr_readdata
	wire   [1:0] mm_interconnect_0_block_dma_csr_address;                     // mm_interconnect_0:block_dma_csr_address -> block_dma:avs_csr_address
	wire         mm_interconnect_0_block_dma_csr_write;                       // mm_interconnect_0:block_dma_csr_write -> block_dma:avs_csr_write
	wire  [31:0] mm_interconnect_0_block_dma_csr_writedata;                   // mm_interconnect_0:block_dma_csr_writedata -> block_dma:avs_csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_program_s1_chipselect;                     // mm_interconnect_0:program_s1_chipselect -> program:chipselect
	wire  [31:0] mm_interconnect_0_program_s1_readdata;                       // program:readdata -> mm_interconnect_0:program_s1_readdata
	wire  [14:0] mm_interconnect_0_program_s1_address;                        // mm_interconnect_0:program_s1_address -> program:address
	wire   [3:0] mm_interconnect_0_program_s1_byteenable;                     // mm_interconnect_0:program_s1_byteenable -> program:byteenable
	wire         mm_interconnect_0_program_s1_write;                          // mm_interconnect_0:program_s1_write -> program:write
	wire  [31:0] mm_interconnect_0_program_s1_writedata;                      // mm_interconnect_0:program_s1_writedata -> program:writedata
	wire         mm_interconnect_0_program_s1_clken;                          // mm_interconnect_0:program_s1_clken -> program:clken
	wire         mm_interconnect_0_dst_ram_s1_chipselect;                     // mm_interconnect_0:dst_ram_s1_chipselect -> dst_ram:chipselect
	wire  [31:0] mm_interconnect_0_dst_ram_s1_readdata;                       // dst_ram:readdata -> mm_interconnect_0:dst_ram_s1_readdata
	wire   [9:0] mm_interconnect_0_dst_ram_s1_address;                        // mm_interconnect_0:dst_ram_s1_address -> dst_ram:address
	wire   [3:0] mm_interconnect_0_dst_ram_s1_byteenable;                     // mm_interconnect_0:dst_ram_s1_byteenable -> dst_ram:byteenable
	wire         mm_interconnect_0_dst_ram_s1_write;                          // mm_interconnect_0:dst_ram_s1_write -> dst_ram:write
	wire  [31:0] mm_interconnect_0_dst_ram_s1_writedata;                      // mm_interconnect_0:dst_ram_s1_writedata -> dst_ram:writedata
	wire         mm_interconnect_0_dst_ram_s1_clken;                          // mm_interconnect_0:dst_ram_s1_clken -> dst_ram:clken
	wire         mm_interconnect_0_src_ram_s1_chipselect;                     // mm_interconnect_0:src_ram_s1_chipselect -> src_ram:chipselect
	wire  [31:0] mm_interconnect_0_src_ram_s1_readdata;                       // src_ram:readdata -> mm_interconnect_0:src_ram_s1_readdata
	wire   [9:0] mm_interconnect_0_src_ram_s1_address;                        // mm_interconnect_0:src_ram_s1_address -> src_ram:address
	wire   [3:0] mm_interconnect_0_src_ram_s1_byteenable;                     // mm_interconnect_0:src_ram_s1_byteenable -> src_ram:byteenable
	wire         mm_interconnect_0_src_ram_s1_write;                          // mm_interconnect_0:src_ram_s1_write -> src_ram:write
	wire  [31:0] mm_interconnect_0_src_ram_s1_writedata;                      // mm_interconnect_0:src_ram_s1_writedata -> src_ram:writedata
	wire         mm_interconnect_0_src_ram_s1_clken;                          // mm_interconnect_0:src_ram_s1_clken -> src_ram:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [block_dma:csi_clock_reset, burst_dma:csi_clock_reset, dst_ram:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, pipelined_dma:csi_clock_reset, program:reset, rst_translator:in_reset, simple_dma:csi_clock_reset, src_ram:reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [dst_ram:reset_req, nios2_gen2_0:reset_req, program:reset_req, rst_translator:reset_req_in, src_ram:reset_req]

	block_transaction_example block_dma (
		.csi_clock_clk                (clk_clk),                                   //        clock.clk
		.csi_clock_reset              (rst_controller_reset_out_reset),            //  clock_reset.reset
		.avm_read_master_read         (block_dma_read_master_read),                //  read_master.read
		.avm_read_master_address      (block_dma_read_master_address),             //             .address
		.avm_read_master_readdata     (block_dma_read_master_readdata),            //             .readdata
		.avm_read_master_waitrequest  (block_dma_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write       (block_dma_write_master_write),              // write_master.write
		.avm_write_master_address     (block_dma_write_master_address),            //             .address
		.avm_write_master_writedata   (block_dma_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest (block_dma_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address              (mm_interconnect_0_block_dma_csr_address),   //          csr.address
		.avs_csr_readdata             (mm_interconnect_0_block_dma_csr_readdata),  //             .readdata
		.avs_csr_write                (mm_interconnect_0_block_dma_csr_write),     //             .write
		.avs_csr_writedata            (mm_interconnect_0_block_dma_csr_writedata)  //             .writedata
	);

	burst_example burst_dma (
		.csi_clock_clk                 (clk_clk),                                   //        clock.clk
		.csi_clock_reset               (rst_controller_reset_out_reset),            //  clock_reset.reset
		.avm_read_master_read          (burst_dma_read_master_read),                //  read_master.read
		.avm_read_master_address       (burst_dma_read_master_address),             //             .address
		.avm_read_master_burstcount    (burst_dma_read_master_burstcount),          //             .burstcount
		.avm_read_master_readdata      (burst_dma_read_master_readdata),            //             .readdata
		.avm_read_master_readdatavalid (burst_dma_read_master_readdatavalid),       //             .readdatavalid
		.avm_read_master_waitrequest   (burst_dma_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write        (burst_dma_write_master_write),              // write_master.write
		.avm_write_master_address      (burst_dma_write_master_address),            //             .address
		.avm_write_master_burstcount   (burst_dma_write_master_burstcount),         //             .burstcount
		.avm_write_master_writedata    (burst_dma_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest  (burst_dma_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address               (mm_interconnect_0_burst_dma_csr_address),   //          csr.address
		.avs_csr_readdata              (mm_interconnect_0_burst_dma_csr_readdata),  //             .readdata
		.avs_csr_write                 (mm_interconnect_0_burst_dma_csr_write),     //             .write
		.avs_csr_writedata             (mm_interconnect_0_burst_dma_csr_writedata)  //             .writedata
	);

	nios_custom_dma_dst_ram dst_ram (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_dst_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_dst_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_dst_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_dst_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_dst_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_dst_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_dst_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	nios_custom_dma_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_custom_dma_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	pipelined_read_example pipelined_dma (
		.csi_clock_clk                 (clk_clk),                                       //        clock.clk
		.csi_clock_reset               (rst_controller_reset_out_reset),                //  clock_reset.reset
		.avm_read_master_read          (pipelined_dma_read_master_read),                //  read_master.read
		.avm_read_master_address       (pipelined_dma_read_master_address),             //             .address
		.avm_read_master_readdata      (pipelined_dma_read_master_readdata),            //             .readdata
		.avm_read_master_readdatavalid (pipelined_dma_read_master_readdatavalid),       //             .readdatavalid
		.avm_read_master_waitrequest   (pipelined_dma_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write        (pipelined_dma_write_master_write),              // write_master.write
		.avm_write_master_address      (pipelined_dma_write_master_address),            //             .address
		.avm_write_master_writedata    (pipelined_dma_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest  (pipelined_dma_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address               (mm_interconnect_0_pipelined_dma_csr_address),   //          csr.address
		.avs_csr_readdata              (mm_interconnect_0_pipelined_dma_csr_readdata),  //             .readdata
		.avs_csr_write                 (mm_interconnect_0_pipelined_dma_csr_write),     //             .write
		.avs_csr_writedata             (mm_interconnect_0_pipelined_dma_csr_writedata)  //             .writedata
	);

	nios_custom_dma_program program_inst (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_program_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_program_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_program_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_program_s1_write),      //       .write
		.readdata   (mm_interconnect_0_program_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_program_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_program_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	simple_example simple_dma (
		.csi_clock_clk                (clk_clk),                                    //        clock.clk
		.csi_clock_reset              (rst_controller_reset_out_reset),             //  clock_reset.reset
		.avm_read_master_read         (simple_dma_read_master_read),                //  read_master.read
		.avm_read_master_address      (simple_dma_read_master_address),             //             .address
		.avm_read_master_readdata     (simple_dma_read_master_readdata),            //             .readdata
		.avm_read_master_waitrequest  (simple_dma_read_master_waitrequest),         //             .waitrequest
		.avm_write_master_write       (simple_dma_write_master_write),              // write_master.write
		.avm_write_master_address     (simple_dma_write_master_address),            //             .address
		.avm_write_master_writedata   (simple_dma_write_master_writedata),          //             .writedata
		.avm_write_master_waitrequest (simple_dma_write_master_waitrequest),        //             .waitrequest
		.avs_csr_address              (mm_interconnect_0_simple_dma_csr_address),   //          csr.address
		.avs_csr_readdata             (mm_interconnect_0_simple_dma_csr_readdata),  //             .readdata
		.avs_csr_write                (mm_interconnect_0_simple_dma_csr_write),     //             .write
		.avs_csr_writedata            (mm_interconnect_0_simple_dma_csr_writedata)  //             .writedata
	);

	nios_custom_dma_src_ram src_ram (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_src_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_src_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_src_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_src_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_src_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_src_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_src_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	nios_custom_dma_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.block_dma_read_master_address                  (block_dma_read_master_address),                               //                    block_dma_read_master.address
		.block_dma_read_master_waitrequest              (block_dma_read_master_waitrequest),                           //                                         .waitrequest
		.block_dma_read_master_read                     (block_dma_read_master_read),                                  //                                         .read
		.block_dma_read_master_readdata                 (block_dma_read_master_readdata),                              //                                         .readdata
		.block_dma_write_master_address                 (block_dma_write_master_address),                              //                   block_dma_write_master.address
		.block_dma_write_master_waitrequest             (block_dma_write_master_waitrequest),                          //                                         .waitrequest
		.block_dma_write_master_write                   (block_dma_write_master_write),                                //                                         .write
		.block_dma_write_master_writedata               (block_dma_write_master_writedata),                            //                                         .writedata
		.burst_dma_read_master_address                  (burst_dma_read_master_address),                               //                    burst_dma_read_master.address
		.burst_dma_read_master_waitrequest              (burst_dma_read_master_waitrequest),                           //                                         .waitrequest
		.burst_dma_read_master_burstcount               (burst_dma_read_master_burstcount),                            //                                         .burstcount
		.burst_dma_read_master_read                     (burst_dma_read_master_read),                                  //                                         .read
		.burst_dma_read_master_readdata                 (burst_dma_read_master_readdata),                              //                                         .readdata
		.burst_dma_read_master_readdatavalid            (burst_dma_read_master_readdatavalid),                         //                                         .readdatavalid
		.burst_dma_write_master_address                 (burst_dma_write_master_address),                              //                   burst_dma_write_master.address
		.burst_dma_write_master_waitrequest             (burst_dma_write_master_waitrequest),                          //                                         .waitrequest
		.burst_dma_write_master_burstcount              (burst_dma_write_master_burstcount),                           //                                         .burstcount
		.burst_dma_write_master_write                   (burst_dma_write_master_write),                                //                                         .write
		.burst_dma_write_master_writedata               (burst_dma_write_master_writedata),                            //                                         .writedata
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.pipelined_dma_read_master_address              (pipelined_dma_read_master_address),                           //                pipelined_dma_read_master.address
		.pipelined_dma_read_master_waitrequest          (pipelined_dma_read_master_waitrequest),                       //                                         .waitrequest
		.pipelined_dma_read_master_read                 (pipelined_dma_read_master_read),                              //                                         .read
		.pipelined_dma_read_master_readdata             (pipelined_dma_read_master_readdata),                          //                                         .readdata
		.pipelined_dma_read_master_readdatavalid        (pipelined_dma_read_master_readdatavalid),                     //                                         .readdatavalid
		.pipelined_dma_write_master_address             (pipelined_dma_write_master_address),                          //               pipelined_dma_write_master.address
		.pipelined_dma_write_master_waitrequest         (pipelined_dma_write_master_waitrequest),                      //                                         .waitrequest
		.pipelined_dma_write_master_write               (pipelined_dma_write_master_write),                            //                                         .write
		.pipelined_dma_write_master_writedata           (pipelined_dma_write_master_writedata),                        //                                         .writedata
		.simple_dma_read_master_address                 (simple_dma_read_master_address),                              //                   simple_dma_read_master.address
		.simple_dma_read_master_waitrequest             (simple_dma_read_master_waitrequest),                          //                                         .waitrequest
		.simple_dma_read_master_read                    (simple_dma_read_master_read),                                 //                                         .read
		.simple_dma_read_master_readdata                (simple_dma_read_master_readdata),                             //                                         .readdata
		.simple_dma_write_master_address                (simple_dma_write_master_address),                             //                  simple_dma_write_master.address
		.simple_dma_write_master_waitrequest            (simple_dma_write_master_waitrequest),                         //                                         .waitrequest
		.simple_dma_write_master_write                  (simple_dma_write_master_write),                               //                                         .write
		.simple_dma_write_master_writedata              (simple_dma_write_master_writedata),                           //                                         .writedata
		.block_dma_csr_address                          (mm_interconnect_0_block_dma_csr_address),                     //                            block_dma_csr.address
		.block_dma_csr_write                            (mm_interconnect_0_block_dma_csr_write),                       //                                         .write
		.block_dma_csr_readdata                         (mm_interconnect_0_block_dma_csr_readdata),                    //                                         .readdata
		.block_dma_csr_writedata                        (mm_interconnect_0_block_dma_csr_writedata),                   //                                         .writedata
		.burst_dma_csr_address                          (mm_interconnect_0_burst_dma_csr_address),                     //                            burst_dma_csr.address
		.burst_dma_csr_write                            (mm_interconnect_0_burst_dma_csr_write),                       //                                         .write
		.burst_dma_csr_readdata                         (mm_interconnect_0_burst_dma_csr_readdata),                    //                                         .readdata
		.burst_dma_csr_writedata                        (mm_interconnect_0_burst_dma_csr_writedata),                   //                                         .writedata
		.dst_ram_s1_address                             (mm_interconnect_0_dst_ram_s1_address),                        //                               dst_ram_s1.address
		.dst_ram_s1_write                               (mm_interconnect_0_dst_ram_s1_write),                          //                                         .write
		.dst_ram_s1_readdata                            (mm_interconnect_0_dst_ram_s1_readdata),                       //                                         .readdata
		.dst_ram_s1_writedata                           (mm_interconnect_0_dst_ram_s1_writedata),                      //                                         .writedata
		.dst_ram_s1_byteenable                          (mm_interconnect_0_dst_ram_s1_byteenable),                     //                                         .byteenable
		.dst_ram_s1_chipselect                          (mm_interconnect_0_dst_ram_s1_chipselect),                     //                                         .chipselect
		.dst_ram_s1_clken                               (mm_interconnect_0_dst_ram_s1_clken),                          //                                         .clken
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.pipelined_dma_csr_address                      (mm_interconnect_0_pipelined_dma_csr_address),                 //                        pipelined_dma_csr.address
		.pipelined_dma_csr_write                        (mm_interconnect_0_pipelined_dma_csr_write),                   //                                         .write
		.pipelined_dma_csr_readdata                     (mm_interconnect_0_pipelined_dma_csr_readdata),                //                                         .readdata
		.pipelined_dma_csr_writedata                    (mm_interconnect_0_pipelined_dma_csr_writedata),               //                                         .writedata
		.program_s1_address                             (mm_interconnect_0_program_s1_address),                        //                               program_s1.address
		.program_s1_write                               (mm_interconnect_0_program_s1_write),                          //                                         .write
		.program_s1_readdata                            (mm_interconnect_0_program_s1_readdata),                       //                                         .readdata
		.program_s1_writedata                           (mm_interconnect_0_program_s1_writedata),                      //                                         .writedata
		.program_s1_byteenable                          (mm_interconnect_0_program_s1_byteenable),                     //                                         .byteenable
		.program_s1_chipselect                          (mm_interconnect_0_program_s1_chipselect),                     //                                         .chipselect
		.program_s1_clken                               (mm_interconnect_0_program_s1_clken),                          //                                         .clken
		.simple_dma_csr_address                         (mm_interconnect_0_simple_dma_csr_address),                    //                           simple_dma_csr.address
		.simple_dma_csr_write                           (mm_interconnect_0_simple_dma_csr_write),                      //                                         .write
		.simple_dma_csr_readdata                        (mm_interconnect_0_simple_dma_csr_readdata),                   //                                         .readdata
		.simple_dma_csr_writedata                       (mm_interconnect_0_simple_dma_csr_writedata),                  //                                         .writedata
		.src_ram_s1_address                             (mm_interconnect_0_src_ram_s1_address),                        //                               src_ram_s1.address
		.src_ram_s1_write                               (mm_interconnect_0_src_ram_s1_write),                          //                                         .write
		.src_ram_s1_readdata                            (mm_interconnect_0_src_ram_s1_readdata),                       //                                         .readdata
		.src_ram_s1_writedata                           (mm_interconnect_0_src_ram_s1_writedata),                      //                                         .writedata
		.src_ram_s1_byteenable                          (mm_interconnect_0_src_ram_s1_byteenable),                     //                                         .byteenable
		.src_ram_s1_chipselect                          (mm_interconnect_0_src_ram_s1_chipselect),                     //                                         .chipselect
		.src_ram_s1_clken                               (mm_interconnect_0_src_ram_s1_clken)                           //                                         .clken
	);

	nios_custom_dma_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
