// dma.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module dma (
		input  wire  clk_clk  // clk.clk
	);

	wire          data_source_pattern_out_valid;                               // data_source:aso_valid -> msgdma_0:st_sink_valid
	wire   [31:0] data_source_pattern_out_data;                                // data_source:aso_data -> msgdma_0:st_sink_data
	wire          data_source_pattern_out_ready;                               // msgdma_0:st_sink_ready -> data_source:aso_ready
	wire          nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire   [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire          nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire          nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire   [17:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire    [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire          nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire          nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire          nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire   [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire          msgdma_0_mm_write_waitrequest;                               // mm_interconnect_0:msgdma_0_mm_write_waitrequest -> msgdma_0:mm_write_waitrequest
	wire   [11:0] msgdma_0_mm_write_address;                                   // msgdma_0:mm_write_address -> mm_interconnect_0:msgdma_0_mm_write_address
	wire    [3:0] msgdma_0_mm_write_byteenable;                                // msgdma_0:mm_write_byteenable -> mm_interconnect_0:msgdma_0_mm_write_byteenable
	wire          msgdma_0_mm_write_write;                                     // msgdma_0:mm_write_write -> mm_interconnect_0:msgdma_0_mm_write_write
	wire   [31:0] msgdma_0_mm_write_writedata;                                 // msgdma_0:mm_write_writedata -> mm_interconnect_0:msgdma_0_mm_write_writedata
	wire   [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire          nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire   [17:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire          nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire          nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire          mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [31:0] mm_interconnect_0_msgdma_0_csr_readdata;                     // msgdma_0:csr_readdata -> mm_interconnect_0:msgdma_0_csr_readdata
	wire    [2:0] mm_interconnect_0_msgdma_0_csr_address;                      // mm_interconnect_0:msgdma_0_csr_address -> msgdma_0:csr_address
	wire          mm_interconnect_0_msgdma_0_csr_read;                         // mm_interconnect_0:msgdma_0_csr_read -> msgdma_0:csr_read
	wire    [3:0] mm_interconnect_0_msgdma_0_csr_byteenable;                   // mm_interconnect_0:msgdma_0_csr_byteenable -> msgdma_0:csr_byteenable
	wire          mm_interconnect_0_msgdma_0_csr_write;                        // mm_interconnect_0:msgdma_0_csr_write -> msgdma_0:csr_write
	wire   [31:0] mm_interconnect_0_msgdma_0_csr_writedata;                    // mm_interconnect_0:msgdma_0_csr_writedata -> msgdma_0:csr_writedata
	wire   [31:0] mm_interconnect_0_data_source_csr_slave_readdata;            // data_source:csr_slave_readdata -> mm_interconnect_0:data_source_csr_slave_readdata
	wire    [2:0] mm_interconnect_0_data_source_csr_slave_address;             // mm_interconnect_0:data_source_csr_slave_address -> data_source:csr_slave_address
	wire          mm_interconnect_0_data_source_csr_slave_read;                // mm_interconnect_0:data_source_csr_slave_read -> data_source:csr_slave_read
	wire    [3:0] mm_interconnect_0_data_source_csr_slave_byteenable;          // mm_interconnect_0:data_source_csr_slave_byteenable -> data_source:csr_slave_byteenable
	wire          mm_interconnect_0_data_source_csr_slave_write;               // mm_interconnect_0:data_source_csr_slave_write -> data_source:csr_slave_write
	wire   [31:0] mm_interconnect_0_data_source_csr_slave_writedata;           // mm_interconnect_0:data_source_csr_slave_writedata -> data_source:csr_slave_writedata
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire          mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest;     // msgdma_0:descriptor_slave_waitrequest -> mm_interconnect_0:msgdma_0_descriptor_slave_waitrequest
	wire   [15:0] mm_interconnect_0_msgdma_0_descriptor_slave_byteenable;      // mm_interconnect_0:msgdma_0_descriptor_slave_byteenable -> msgdma_0:descriptor_slave_byteenable
	wire          mm_interconnect_0_msgdma_0_descriptor_slave_write;           // mm_interconnect_0:msgdma_0_descriptor_slave_write -> msgdma_0:descriptor_slave_write
	wire  [127:0] mm_interconnect_0_msgdma_0_descriptor_slave_writedata;       // mm_interconnect_0:msgdma_0_descriptor_slave_writedata -> msgdma_0:descriptor_slave_writedata
	wire          mm_interconnect_0_ocram_s1_chipselect;                       // mm_interconnect_0:ocram_s1_chipselect -> ocram:chipselect
	wire   [31:0] mm_interconnect_0_ocram_s1_readdata;                         // ocram:readdata -> mm_interconnect_0:ocram_s1_readdata
	wire   [13:0] mm_interconnect_0_ocram_s1_address;                          // mm_interconnect_0:ocram_s1_address -> ocram:address
	wire    [3:0] mm_interconnect_0_ocram_s1_byteenable;                       // mm_interconnect_0:ocram_s1_byteenable -> ocram:byteenable
	wire          mm_interconnect_0_ocram_s1_write;                            // mm_interconnect_0:ocram_s1_write -> ocram:write
	wire   [31:0] mm_interconnect_0_ocram_s1_writedata;                        // mm_interconnect_0:ocram_s1_writedata -> ocram:writedata
	wire          mm_interconnect_0_ocram_s1_clken;                            // mm_interconnect_0:ocram_s1_clken -> ocram:clken
	wire          mm_interconnect_0_data_destination_s1_chipselect;            // mm_interconnect_0:data_destination_s1_chipselect -> data_destination:chipselect
	wire   [31:0] mm_interconnect_0_data_destination_s1_readdata;              // data_destination:readdata -> mm_interconnect_0:data_destination_s1_readdata
	wire    [9:0] mm_interconnect_0_data_destination_s1_address;               // mm_interconnect_0:data_destination_s1_address -> data_destination:address
	wire    [3:0] mm_interconnect_0_data_destination_s1_byteenable;            // mm_interconnect_0:data_destination_s1_byteenable -> data_destination:byteenable
	wire          mm_interconnect_0_data_destination_s1_write;                 // mm_interconnect_0:data_destination_s1_write -> data_destination:write
	wire   [31:0] mm_interconnect_0_data_destination_s1_writedata;             // mm_interconnect_0:data_destination_s1_writedata -> data_destination:writedata
	wire          mm_interconnect_0_data_destination_s1_clken;                 // mm_interconnect_0:data_destination_s1_clken -> data_destination:clken
	wire          irq_mapper_receiver0_irq;                                    // msgdma_0:csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire   [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire          rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [data_destination:reset, data_source:reset_reset, mm_interconnect_0:msgdma_0_reset_n_reset_bridge_in_reset_reset, msgdma_0:reset_n_reset_n, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [data_destination:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, ocram:reset, rst_translator_001:in_reset]
	wire          rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, ocram:reset_req, rst_translator_001:reset_req_in]

	dma_data_destination data_destination (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_data_destination_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_destination_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_destination_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_destination_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_destination_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_destination_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_destination_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	dma_data_source #(
		.ST_DATA_W            (32),
		.BYPASS_ENABLED       (0),
		.AVALON_ENABLED       (1),
		.CROSS_CLK_SYNC_DEPTH (2)
	) data_source (
		.csr_clk_clk          (clk_clk),                                            //         csr_clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                     //           reset.reset
		.csr_slave_address    (mm_interconnect_0_data_source_csr_slave_address),    //       csr_slave.address
		.csr_slave_write      (mm_interconnect_0_data_source_csr_slave_write),      //                .write
		.csr_slave_read       (mm_interconnect_0_data_source_csr_slave_read),       //                .read
		.csr_slave_byteenable (mm_interconnect_0_data_source_csr_slave_byteenable), //                .byteenable
		.csr_slave_writedata  (mm_interconnect_0_data_source_csr_slave_writedata),  //                .writedata
		.csr_slave_readdata   (mm_interconnect_0_data_source_csr_slave_readdata),   //                .readdata
		.pattern_out_clk_clk  (clk_clk),                                            // pattern_out_clk.clk
		.aso_valid            (data_source_pattern_out_valid),                      //     pattern_out.valid
		.aso_ready            (data_source_pattern_out_ready),                      //                .ready
		.aso_data             (data_source_pattern_out_data)                        //                .data
	);

	dma_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	dma_msgdma_0 msgdma_0 (
		.mm_write_address             (msgdma_0_mm_write_address),                               //         mm_write.address
		.mm_write_write               (msgdma_0_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (msgdma_0_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (msgdma_0_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (msgdma_0_mm_write_waitrequest),                           //                 .waitrequest
		.clock_clk                    (clk_clk),                                                 //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                         //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_msgdma_0_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_msgdma_0_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_msgdma_0_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_msgdma_0_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_msgdma_0_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_msgdma_0_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_msgdma_0_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_msgdma_0_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_msgdma_0_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver0_irq),                                //          csr_irq.irq
		.st_sink_data                 (data_source_pattern_out_data),                            //          st_sink.data
		.st_sink_valid                (data_source_pattern_out_valid),                           //                 .valid
		.st_sink_ready                (data_source_pattern_out_ready)                            //                 .ready
	);

	dma_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	dma_ocram ocram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ocram_s1_address),     //     s1.address
		.clken      (mm_interconnect_0_ocram_s1_clken),       //       .clken
		.chipselect (mm_interconnect_0_ocram_s1_chipselect),  //       .chipselect
		.write      (mm_interconnect_0_ocram_s1_write),       //       .write
		.readdata   (mm_interconnect_0_ocram_s1_readdata),    //       .readdata
		.writedata  (mm_interconnect_0_ocram_s1_writedata),   //       .writedata
		.byteenable (mm_interconnect_0_ocram_s1_byteenable),  //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	dma_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.msgdma_0_reset_n_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                              //   msgdma_0_reset_n_reset_bridge_in_reset.reset
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.msgdma_0_mm_write_address                      (msgdma_0_mm_write_address),                                   //                        msgdma_0_mm_write.address
		.msgdma_0_mm_write_waitrequest                  (msgdma_0_mm_write_waitrequest),                               //                                         .waitrequest
		.msgdma_0_mm_write_byteenable                   (msgdma_0_mm_write_byteenable),                                //                                         .byteenable
		.msgdma_0_mm_write_write                        (msgdma_0_mm_write_write),                                     //                                         .write
		.msgdma_0_mm_write_writedata                    (msgdma_0_mm_write_writedata),                                 //                                         .writedata
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.data_destination_s1_address                    (mm_interconnect_0_data_destination_s1_address),               //                      data_destination_s1.address
		.data_destination_s1_write                      (mm_interconnect_0_data_destination_s1_write),                 //                                         .write
		.data_destination_s1_readdata                   (mm_interconnect_0_data_destination_s1_readdata),              //                                         .readdata
		.data_destination_s1_writedata                  (mm_interconnect_0_data_destination_s1_writedata),             //                                         .writedata
		.data_destination_s1_byteenable                 (mm_interconnect_0_data_destination_s1_byteenable),            //                                         .byteenable
		.data_destination_s1_chipselect                 (mm_interconnect_0_data_destination_s1_chipselect),            //                                         .chipselect
		.data_destination_s1_clken                      (mm_interconnect_0_data_destination_s1_clken),                 //                                         .clken
		.data_source_csr_slave_address                  (mm_interconnect_0_data_source_csr_slave_address),             //                    data_source_csr_slave.address
		.data_source_csr_slave_write                    (mm_interconnect_0_data_source_csr_slave_write),               //                                         .write
		.data_source_csr_slave_read                     (mm_interconnect_0_data_source_csr_slave_read),                //                                         .read
		.data_source_csr_slave_readdata                 (mm_interconnect_0_data_source_csr_slave_readdata),            //                                         .readdata
		.data_source_csr_slave_writedata                (mm_interconnect_0_data_source_csr_slave_writedata),           //                                         .writedata
		.data_source_csr_slave_byteenable               (mm_interconnect_0_data_source_csr_slave_byteenable),          //                                         .byteenable
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.msgdma_0_csr_address                           (mm_interconnect_0_msgdma_0_csr_address),                      //                             msgdma_0_csr.address
		.msgdma_0_csr_write                             (mm_interconnect_0_msgdma_0_csr_write),                        //                                         .write
		.msgdma_0_csr_read                              (mm_interconnect_0_msgdma_0_csr_read),                         //                                         .read
		.msgdma_0_csr_readdata                          (mm_interconnect_0_msgdma_0_csr_readdata),                     //                                         .readdata
		.msgdma_0_csr_writedata                         (mm_interconnect_0_msgdma_0_csr_writedata),                    //                                         .writedata
		.msgdma_0_csr_byteenable                        (mm_interconnect_0_msgdma_0_csr_byteenable),                   //                                         .byteenable
		.msgdma_0_descriptor_slave_write                (mm_interconnect_0_msgdma_0_descriptor_slave_write),           //                msgdma_0_descriptor_slave.write
		.msgdma_0_descriptor_slave_writedata            (mm_interconnect_0_msgdma_0_descriptor_slave_writedata),       //                                         .writedata
		.msgdma_0_descriptor_slave_byteenable           (mm_interconnect_0_msgdma_0_descriptor_slave_byteenable),      //                                         .byteenable
		.msgdma_0_descriptor_slave_waitrequest          (mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest),     //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.ocram_s1_address                               (mm_interconnect_0_ocram_s1_address),                          //                                 ocram_s1.address
		.ocram_s1_write                                 (mm_interconnect_0_ocram_s1_write),                            //                                         .write
		.ocram_s1_readdata                              (mm_interconnect_0_ocram_s1_readdata),                         //                                         .readdata
		.ocram_s1_writedata                             (mm_interconnect_0_ocram_s1_writedata),                        //                                         .writedata
		.ocram_s1_byteenable                            (mm_interconnect_0_ocram_s1_byteenable),                       //                                         .byteenable
		.ocram_s1_chipselect                            (mm_interconnect_0_ocram_s1_chipselect),                       //                                         .chipselect
		.ocram_s1_clken                                 (mm_interconnect_0_ocram_s1_clken)                             //                                         .clken
	);

	dma_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
