// HelloNiosIntr.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module HelloNiosIntr (
		input  wire  clk_clk  // clk.clk
	);

	wire         niosintr_debug_reset_request_reset;                     // NiosIntr:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] niosintr_data_master_readdata;                          // mm_interconnect_0:NiosIntr_data_master_readdata -> NiosIntr:d_readdata
	wire         niosintr_data_master_waitrequest;                       // mm_interconnect_0:NiosIntr_data_master_waitrequest -> NiosIntr:d_waitrequest
	wire         niosintr_data_master_debugaccess;                       // NiosIntr:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosIntr_data_master_debugaccess
	wire  [17:0] niosintr_data_master_address;                           // NiosIntr:d_address -> mm_interconnect_0:NiosIntr_data_master_address
	wire   [3:0] niosintr_data_master_byteenable;                        // NiosIntr:d_byteenable -> mm_interconnect_0:NiosIntr_data_master_byteenable
	wire         niosintr_data_master_read;                              // NiosIntr:d_read -> mm_interconnect_0:NiosIntr_data_master_read
	wire         niosintr_data_master_readdatavalid;                     // mm_interconnect_0:NiosIntr_data_master_readdatavalid -> NiosIntr:d_readdatavalid
	wire         niosintr_data_master_write;                             // NiosIntr:d_write -> mm_interconnect_0:NiosIntr_data_master_write
	wire  [31:0] niosintr_data_master_writedata;                         // NiosIntr:d_writedata -> mm_interconnect_0:NiosIntr_data_master_writedata
	wire  [31:0] niosintr_instruction_master_readdata;                   // mm_interconnect_0:NiosIntr_instruction_master_readdata -> NiosIntr:i_readdata
	wire         niosintr_instruction_master_waitrequest;                // mm_interconnect_0:NiosIntr_instruction_master_waitrequest -> NiosIntr:i_waitrequest
	wire  [17:0] niosintr_instruction_master_address;                    // NiosIntr:i_address -> mm_interconnect_0:NiosIntr_instruction_master_address
	wire         niosintr_instruction_master_read;                       // NiosIntr:i_read -> mm_interconnect_0:NiosIntr_instruction_master_read
	wire         niosintr_instruction_master_readdatavalid;              // mm_interconnect_0:NiosIntr_instruction_master_readdatavalid -> NiosIntr:i_readdatavalid
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;     // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;  // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;      // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;         // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;    // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_niosintr_debug_mem_slave_readdata;    // NiosIntr:debug_mem_slave_readdata -> mm_interconnect_0:NiosIntr_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosintr_debug_mem_slave_waitrequest; // NiosIntr:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosIntr_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosintr_debug_mem_slave_debugaccess; // mm_interconnect_0:NiosIntr_debug_mem_slave_debugaccess -> NiosIntr:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosintr_debug_mem_slave_address;     // mm_interconnect_0:NiosIntr_debug_mem_slave_address -> NiosIntr:debug_mem_slave_address
	wire         mm_interconnect_0_niosintr_debug_mem_slave_read;        // mm_interconnect_0:NiosIntr_debug_mem_slave_read -> NiosIntr:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosintr_debug_mem_slave_byteenable;  // mm_interconnect_0:NiosIntr_debug_mem_slave_byteenable -> NiosIntr:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosintr_debug_mem_slave_write;       // mm_interconnect_0:NiosIntr_debug_mem_slave_write -> NiosIntr:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosintr_debug_mem_slave_writedata;   // mm_interconnect_0:NiosIntr_debug_mem_slave_writedata -> NiosIntr:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                   // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                     // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [13:0] mm_interconnect_0_sram_s1_address;                      // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                   // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                        // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                    // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                        // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                  // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                    // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                     // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                       // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                   // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         irq_mapper_receiver0_irq;                               // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                               // TIMER:irq -> irq_mapper:receiver1_irq
	wire  [31:0] niosintr_irq_irq;                                       // irq_mapper:sender_irq -> NiosIntr:irq
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [DEBUG:rst_n, NiosIntr:reset_n, SRAM:reset, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:NiosIntr_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [NiosIntr:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	HelloNiosIntr_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	HelloNiosIntr_NiosIntr niosintr (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (niosintr_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosintr_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosintr_data_master_read),                              //                          .read
		.d_readdata                          (niosintr_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosintr_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosintr_data_master_write),                             //                          .write
		.d_writedata                         (niosintr_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (niosintr_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (niosintr_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosintr_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosintr_instruction_master_read),                       //                          .read
		.i_readdata                          (niosintr_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosintr_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (niosintr_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosintr_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosintr_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosintr_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosintr_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosintr_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosintr_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosintr_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosintr_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosintr_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosintr_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	HelloNiosIntr_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	HelloNiosIntr_TIMER timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	HelloNiosIntr_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                              (clk_clk),                                                //                            clk_0_clk.clk
		.NiosIntr_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                         // NiosIntr_reset_reset_bridge_in_reset.reset
		.NiosIntr_data_master_address               (niosintr_data_master_address),                           //                 NiosIntr_data_master.address
		.NiosIntr_data_master_waitrequest           (niosintr_data_master_waitrequest),                       //                                     .waitrequest
		.NiosIntr_data_master_byteenable            (niosintr_data_master_byteenable),                        //                                     .byteenable
		.NiosIntr_data_master_read                  (niosintr_data_master_read),                              //                                     .read
		.NiosIntr_data_master_readdata              (niosintr_data_master_readdata),                          //                                     .readdata
		.NiosIntr_data_master_readdatavalid         (niosintr_data_master_readdatavalid),                     //                                     .readdatavalid
		.NiosIntr_data_master_write                 (niosintr_data_master_write),                             //                                     .write
		.NiosIntr_data_master_writedata             (niosintr_data_master_writedata),                         //                                     .writedata
		.NiosIntr_data_master_debugaccess           (niosintr_data_master_debugaccess),                       //                                     .debugaccess
		.NiosIntr_instruction_master_address        (niosintr_instruction_master_address),                    //          NiosIntr_instruction_master.address
		.NiosIntr_instruction_master_waitrequest    (niosintr_instruction_master_waitrequest),                //                                     .waitrequest
		.NiosIntr_instruction_master_read           (niosintr_instruction_master_read),                       //                                     .read
		.NiosIntr_instruction_master_readdata       (niosintr_instruction_master_readdata),                   //                                     .readdata
		.NiosIntr_instruction_master_readdatavalid  (niosintr_instruction_master_readdatavalid),              //                                     .readdatavalid
		.DEBUG_avalon_jtag_slave_address            (mm_interconnect_0_debug_avalon_jtag_slave_address),      //              DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write              (mm_interconnect_0_debug_avalon_jtag_slave_write),        //                                     .write
		.DEBUG_avalon_jtag_slave_read               (mm_interconnect_0_debug_avalon_jtag_slave_read),         //                                     .read
		.DEBUG_avalon_jtag_slave_readdata           (mm_interconnect_0_debug_avalon_jtag_slave_readdata),     //                                     .readdata
		.DEBUG_avalon_jtag_slave_writedata          (mm_interconnect_0_debug_avalon_jtag_slave_writedata),    //                                     .writedata
		.DEBUG_avalon_jtag_slave_waitrequest        (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),  //                                     .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect         (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),   //                                     .chipselect
		.NiosIntr_debug_mem_slave_address           (mm_interconnect_0_niosintr_debug_mem_slave_address),     //             NiosIntr_debug_mem_slave.address
		.NiosIntr_debug_mem_slave_write             (mm_interconnect_0_niosintr_debug_mem_slave_write),       //                                     .write
		.NiosIntr_debug_mem_slave_read              (mm_interconnect_0_niosintr_debug_mem_slave_read),        //                                     .read
		.NiosIntr_debug_mem_slave_readdata          (mm_interconnect_0_niosintr_debug_mem_slave_readdata),    //                                     .readdata
		.NiosIntr_debug_mem_slave_writedata         (mm_interconnect_0_niosintr_debug_mem_slave_writedata),   //                                     .writedata
		.NiosIntr_debug_mem_slave_byteenable        (mm_interconnect_0_niosintr_debug_mem_slave_byteenable),  //                                     .byteenable
		.NiosIntr_debug_mem_slave_waitrequest       (mm_interconnect_0_niosintr_debug_mem_slave_waitrequest), //                                     .waitrequest
		.NiosIntr_debug_mem_slave_debugaccess       (mm_interconnect_0_niosintr_debug_mem_slave_debugaccess), //                                     .debugaccess
		.SRAM_s1_address                            (mm_interconnect_0_sram_s1_address),                      //                              SRAM_s1.address
		.SRAM_s1_write                              (mm_interconnect_0_sram_s1_write),                        //                                     .write
		.SRAM_s1_readdata                           (mm_interconnect_0_sram_s1_readdata),                     //                                     .readdata
		.SRAM_s1_writedata                          (mm_interconnect_0_sram_s1_writedata),                    //                                     .writedata
		.SRAM_s1_byteenable                         (mm_interconnect_0_sram_s1_byteenable),                   //                                     .byteenable
		.SRAM_s1_chipselect                         (mm_interconnect_0_sram_s1_chipselect),                   //                                     .chipselect
		.SRAM_s1_clken                              (mm_interconnect_0_sram_s1_clken),                        //                                     .clken
		.TIMER_s1_address                           (mm_interconnect_0_timer_s1_address),                     //                             TIMER_s1.address
		.TIMER_s1_write                             (mm_interconnect_0_timer_s1_write),                       //                                     .write
		.TIMER_s1_readdata                          (mm_interconnect_0_timer_s1_readdata),                    //                                     .readdata
		.TIMER_s1_writedata                         (mm_interconnect_0_timer_s1_writedata),                   //                                     .writedata
		.TIMER_s1_chipselect                        (mm_interconnect_0_timer_s1_chipselect)                   //                                     .chipselect
	);

	HelloNiosIntr_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (niosintr_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (niosintr_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
