
module NiosInst (
	clk_clk);	

	input		clk_clk;
endmodule
