// Nios_Buffer.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module Nios_Buffer (
		input  wire  clk_clk  // clk.clk
	);

	wire         nios_buff_debug_reset_request_reset;                     // NIOS_BUFF:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nios_buff_data_master_readdata;                          // mm_interconnect_0:NIOS_BUFF_data_master_readdata -> NIOS_BUFF:d_readdata
	wire         nios_buff_data_master_waitrequest;                       // mm_interconnect_0:NIOS_BUFF_data_master_waitrequest -> NIOS_BUFF:d_waitrequest
	wire         nios_buff_data_master_debugaccess;                       // NIOS_BUFF:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS_BUFF_data_master_debugaccess
	wire  [17:0] nios_buff_data_master_address;                           // NIOS_BUFF:d_address -> mm_interconnect_0:NIOS_BUFF_data_master_address
	wire   [3:0] nios_buff_data_master_byteenable;                        // NIOS_BUFF:d_byteenable -> mm_interconnect_0:NIOS_BUFF_data_master_byteenable
	wire         nios_buff_data_master_read;                              // NIOS_BUFF:d_read -> mm_interconnect_0:NIOS_BUFF_data_master_read
	wire         nios_buff_data_master_readdatavalid;                     // mm_interconnect_0:NIOS_BUFF_data_master_readdatavalid -> NIOS_BUFF:d_readdatavalid
	wire         nios_buff_data_master_write;                             // NIOS_BUFF:d_write -> mm_interconnect_0:NIOS_BUFF_data_master_write
	wire  [31:0] nios_buff_data_master_writedata;                         // NIOS_BUFF:d_writedata -> mm_interconnect_0:NIOS_BUFF_data_master_writedata
	wire  [31:0] nios_buff_instruction_master_readdata;                   // mm_interconnect_0:NIOS_BUFF_instruction_master_readdata -> NIOS_BUFF:i_readdata
	wire         nios_buff_instruction_master_waitrequest;                // mm_interconnect_0:NIOS_BUFF_instruction_master_waitrequest -> NIOS_BUFF:i_waitrequest
	wire  [17:0] nios_buff_instruction_master_address;                    // NIOS_BUFF:i_address -> mm_interconnect_0:NIOS_BUFF_instruction_master_address
	wire         nios_buff_instruction_master_read;                       // NIOS_BUFF:i_read -> mm_interconnect_0:NIOS_BUFF_instruction_master_read
	wire         nios_buff_instruction_master_readdatavalid;              // mm_interconnect_0:NIOS_BUFF_instruction_master_readdatavalid -> NIOS_BUFF:i_readdatavalid
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;    // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;      // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;   // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;          // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;         // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire         mm_interconnect_0_mybuffer_avalon_slave_0_chipselect;    // mm_interconnect_0:MyBuffer_avalon_slave_0_chipselect -> MyBuffer:chipselect
	wire  [31:0] mm_interconnect_0_mybuffer_avalon_slave_0_readdata;      // MyBuffer:readdata -> mm_interconnect_0:MyBuffer_avalon_slave_0_readdata
	wire   [9:0] mm_interconnect_0_mybuffer_avalon_slave_0_address;       // mm_interconnect_0:MyBuffer_avalon_slave_0_address -> MyBuffer:address
	wire         mm_interconnect_0_mybuffer_avalon_slave_0_read;          // mm_interconnect_0:MyBuffer_avalon_slave_0_read -> MyBuffer:read
	wire         mm_interconnect_0_mybuffer_avalon_slave_0_write;         // mm_interconnect_0:MyBuffer_avalon_slave_0_write -> MyBuffer:write
	wire  [31:0] mm_interconnect_0_mybuffer_avalon_slave_0_writedata;     // mm_interconnect_0:MyBuffer_avalon_slave_0_writedata -> MyBuffer:writedata
	wire  [31:0] mm_interconnect_0_nios_buff_debug_mem_slave_readdata;    // NIOS_BUFF:debug_mem_slave_readdata -> mm_interconnect_0:NIOS_BUFF_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_buff_debug_mem_slave_waitrequest; // NIOS_BUFF:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS_BUFF_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_buff_debug_mem_slave_debugaccess; // mm_interconnect_0:NIOS_BUFF_debug_mem_slave_debugaccess -> NIOS_BUFF:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_buff_debug_mem_slave_address;     // mm_interconnect_0:NIOS_BUFF_debug_mem_slave_address -> NIOS_BUFF:debug_mem_slave_address
	wire         mm_interconnect_0_nios_buff_debug_mem_slave_read;        // mm_interconnect_0:NIOS_BUFF_debug_mem_slave_read -> NIOS_BUFF:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_buff_debug_mem_slave_byteenable;  // mm_interconnect_0:NIOS_BUFF_debug_mem_slave_byteenable -> NIOS_BUFF:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_buff_debug_mem_slave_write;       // mm_interconnect_0:NIOS_BUFF_debug_mem_slave_write -> NIOS_BUFF:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_buff_debug_mem_slave_writedata;   // mm_interconnect_0:NIOS_BUFF_debug_mem_slave_writedata -> NIOS_BUFF:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                    // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                      // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [13:0] mm_interconnect_0_sram_s1_address;                       // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                    // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                         // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                     // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                         // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         irq_mapper_receiver0_irq;                                // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios_buff_irq_irq;                                       // irq_mapper:sender_irq -> NIOS_BUFF:irq
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [DEBUG:rst_n, MyBuffer:reset_n, NIOS_BUFF:reset_n, SRAM:reset, irq_mapper:reset, mm_interconnect_0:NIOS_BUFF_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                      // rst_controller:reset_req -> [NIOS_BUFF:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	Nios_Buffer_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	CustomIP mybuffer (
		.address    (mm_interconnect_0_mybuffer_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_mybuffer_avalon_slave_0_chipselect), //               .chipselect
		.read       (mm_interconnect_0_mybuffer_avalon_slave_0_read),       //               .read
		.write      (mm_interconnect_0_mybuffer_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_mybuffer_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_mybuffer_avalon_slave_0_readdata),   //               .readdata
		.clk        (clk_clk),                                              //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset)                       //          reset.reset_n
	);

	Nios_Buffer_NIOS_BUFF nios_buff (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (nios_buff_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_buff_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_buff_data_master_read),                              //                          .read
		.d_readdata                          (nios_buff_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_buff_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_buff_data_master_write),                             //                          .write
		.d_writedata                         (nios_buff_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_buff_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_buff_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_buff_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_buff_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_buff_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_buff_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_buff_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_buff_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_buff_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_buff_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_buff_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_buff_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_buff_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_buff_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_buff_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_buff_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_buff_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	Nios_Buffer_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	Nios_Buffer_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                               (clk_clk),                                                 //                             clk_0_clk.clk
		.NIOS_BUFF_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // NIOS_BUFF_reset_reset_bridge_in_reset.reset
		.NIOS_BUFF_data_master_address               (nios_buff_data_master_address),                           //                 NIOS_BUFF_data_master.address
		.NIOS_BUFF_data_master_waitrequest           (nios_buff_data_master_waitrequest),                       //                                      .waitrequest
		.NIOS_BUFF_data_master_byteenable            (nios_buff_data_master_byteenable),                        //                                      .byteenable
		.NIOS_BUFF_data_master_read                  (nios_buff_data_master_read),                              //                                      .read
		.NIOS_BUFF_data_master_readdata              (nios_buff_data_master_readdata),                          //                                      .readdata
		.NIOS_BUFF_data_master_readdatavalid         (nios_buff_data_master_readdatavalid),                     //                                      .readdatavalid
		.NIOS_BUFF_data_master_write                 (nios_buff_data_master_write),                             //                                      .write
		.NIOS_BUFF_data_master_writedata             (nios_buff_data_master_writedata),                         //                                      .writedata
		.NIOS_BUFF_data_master_debugaccess           (nios_buff_data_master_debugaccess),                       //                                      .debugaccess
		.NIOS_BUFF_instruction_master_address        (nios_buff_instruction_master_address),                    //          NIOS_BUFF_instruction_master.address
		.NIOS_BUFF_instruction_master_waitrequest    (nios_buff_instruction_master_waitrequest),                //                                      .waitrequest
		.NIOS_BUFF_instruction_master_read           (nios_buff_instruction_master_read),                       //                                      .read
		.NIOS_BUFF_instruction_master_readdata       (nios_buff_instruction_master_readdata),                   //                                      .readdata
		.NIOS_BUFF_instruction_master_readdatavalid  (nios_buff_instruction_master_readdatavalid),              //                                      .readdatavalid
		.DEBUG_avalon_jtag_slave_address             (mm_interconnect_0_debug_avalon_jtag_slave_address),       //               DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write               (mm_interconnect_0_debug_avalon_jtag_slave_write),         //                                      .write
		.DEBUG_avalon_jtag_slave_read                (mm_interconnect_0_debug_avalon_jtag_slave_read),          //                                      .read
		.DEBUG_avalon_jtag_slave_readdata            (mm_interconnect_0_debug_avalon_jtag_slave_readdata),      //                                      .readdata
		.DEBUG_avalon_jtag_slave_writedata           (mm_interconnect_0_debug_avalon_jtag_slave_writedata),     //                                      .writedata
		.DEBUG_avalon_jtag_slave_waitrequest         (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),   //                                      .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect          (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),    //                                      .chipselect
		.MyBuffer_avalon_slave_0_address             (mm_interconnect_0_mybuffer_avalon_slave_0_address),       //               MyBuffer_avalon_slave_0.address
		.MyBuffer_avalon_slave_0_write               (mm_interconnect_0_mybuffer_avalon_slave_0_write),         //                                      .write
		.MyBuffer_avalon_slave_0_read                (mm_interconnect_0_mybuffer_avalon_slave_0_read),          //                                      .read
		.MyBuffer_avalon_slave_0_readdata            (mm_interconnect_0_mybuffer_avalon_slave_0_readdata),      //                                      .readdata
		.MyBuffer_avalon_slave_0_writedata           (mm_interconnect_0_mybuffer_avalon_slave_0_writedata),     //                                      .writedata
		.MyBuffer_avalon_slave_0_chipselect          (mm_interconnect_0_mybuffer_avalon_slave_0_chipselect),    //                                      .chipselect
		.NIOS_BUFF_debug_mem_slave_address           (mm_interconnect_0_nios_buff_debug_mem_slave_address),     //             NIOS_BUFF_debug_mem_slave.address
		.NIOS_BUFF_debug_mem_slave_write             (mm_interconnect_0_nios_buff_debug_mem_slave_write),       //                                      .write
		.NIOS_BUFF_debug_mem_slave_read              (mm_interconnect_0_nios_buff_debug_mem_slave_read),        //                                      .read
		.NIOS_BUFF_debug_mem_slave_readdata          (mm_interconnect_0_nios_buff_debug_mem_slave_readdata),    //                                      .readdata
		.NIOS_BUFF_debug_mem_slave_writedata         (mm_interconnect_0_nios_buff_debug_mem_slave_writedata),   //                                      .writedata
		.NIOS_BUFF_debug_mem_slave_byteenable        (mm_interconnect_0_nios_buff_debug_mem_slave_byteenable),  //                                      .byteenable
		.NIOS_BUFF_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_buff_debug_mem_slave_waitrequest), //                                      .waitrequest
		.NIOS_BUFF_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_buff_debug_mem_slave_debugaccess), //                                      .debugaccess
		.SRAM_s1_address                             (mm_interconnect_0_sram_s1_address),                       //                               SRAM_s1.address
		.SRAM_s1_write                               (mm_interconnect_0_sram_s1_write),                         //                                      .write
		.SRAM_s1_readdata                            (mm_interconnect_0_sram_s1_readdata),                      //                                      .readdata
		.SRAM_s1_writedata                           (mm_interconnect_0_sram_s1_writedata),                     //                                      .writedata
		.SRAM_s1_byteenable                          (mm_interconnect_0_sram_s1_byteenable),                    //                                      .byteenable
		.SRAM_s1_chipselect                          (mm_interconnect_0_sram_s1_chipselect),                    //                                      .chipselect
		.SRAM_s1_clken                               (mm_interconnect_0_sram_s1_clken)                          //                                      .clken
	);

	Nios_Buffer_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios_buff_irq_irq)               //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios_buff_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
