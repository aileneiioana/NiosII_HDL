// Nios_Custom_IP2.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module Nios_Custom_IP2 (
		input  wire  clk_clk  // clk.clk
	);

	wire         nioscustomip2_debug_reset_request_reset;                     // NiosCustomIP2:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nioscustomip2_data_master_readdata;                          // mm_interconnect_0:NiosCustomIP2_data_master_readdata -> NiosCustomIP2:d_readdata
	wire         nioscustomip2_data_master_waitrequest;                       // mm_interconnect_0:NiosCustomIP2_data_master_waitrequest -> NiosCustomIP2:d_waitrequest
	wire         nioscustomip2_data_master_debugaccess;                       // NiosCustomIP2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosCustomIP2_data_master_debugaccess
	wire  [17:0] nioscustomip2_data_master_address;                           // NiosCustomIP2:d_address -> mm_interconnect_0:NiosCustomIP2_data_master_address
	wire   [3:0] nioscustomip2_data_master_byteenable;                        // NiosCustomIP2:d_byteenable -> mm_interconnect_0:NiosCustomIP2_data_master_byteenable
	wire         nioscustomip2_data_master_read;                              // NiosCustomIP2:d_read -> mm_interconnect_0:NiosCustomIP2_data_master_read
	wire         nioscustomip2_data_master_write;                             // NiosCustomIP2:d_write -> mm_interconnect_0:NiosCustomIP2_data_master_write
	wire  [31:0] nioscustomip2_data_master_writedata;                         // NiosCustomIP2:d_writedata -> mm_interconnect_0:NiosCustomIP2_data_master_writedata
	wire  [31:0] nioscustomip2_instruction_master_readdata;                   // mm_interconnect_0:NiosCustomIP2_instruction_master_readdata -> NiosCustomIP2:i_readdata
	wire         nioscustomip2_instruction_master_waitrequest;                // mm_interconnect_0:NiosCustomIP2_instruction_master_waitrequest -> NiosCustomIP2:i_waitrequest
	wire  [17:0] nioscustomip2_instruction_master_address;                    // NiosCustomIP2:i_address -> mm_interconnect_0:NiosCustomIP2_instruction_master_address
	wire         nioscustomip2_instruction_master_read;                       // NiosCustomIP2:i_read -> mm_interconnect_0:NiosCustomIP2_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;          // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;       // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;           // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;              // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;             // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;         // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire         mm_interconnect_0_myreg_0_avalon_slave_0_chipselect;         // mm_interconnect_0:MyReg_0_avalon_slave_0_chipselect -> MyReg_0:chipselect
	wire  [31:0] mm_interconnect_0_myreg_0_avalon_slave_0_readdata;           // MyReg_0:readdata -> mm_interconnect_0:MyReg_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_myreg_0_avalon_slave_0_address;            // mm_interconnect_0:MyReg_0_avalon_slave_0_address -> MyReg_0:address
	wire         mm_interconnect_0_myreg_0_avalon_slave_0_read;               // mm_interconnect_0:MyReg_0_avalon_slave_0_read -> MyReg_0:read
	wire         mm_interconnect_0_myreg_0_avalon_slave_0_write;              // mm_interconnect_0:MyReg_0_avalon_slave_0_write -> MyReg_0:write
	wire  [31:0] mm_interconnect_0_myreg_0_avalon_slave_0_writedata;          // mm_interconnect_0:MyReg_0_avalon_slave_0_writedata -> MyReg_0:writedata
	wire  [31:0] mm_interconnect_0_nioscustomip2_debug_mem_slave_readdata;    // NiosCustomIP2:debug_mem_slave_readdata -> mm_interconnect_0:NiosCustomIP2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nioscustomip2_debug_mem_slave_waitrequest; // NiosCustomIP2:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosCustomIP2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nioscustomip2_debug_mem_slave_debugaccess; // mm_interconnect_0:NiosCustomIP2_debug_mem_slave_debugaccess -> NiosCustomIP2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nioscustomip2_debug_mem_slave_address;     // mm_interconnect_0:NiosCustomIP2_debug_mem_slave_address -> NiosCustomIP2:debug_mem_slave_address
	wire         mm_interconnect_0_nioscustomip2_debug_mem_slave_read;        // mm_interconnect_0:NiosCustomIP2_debug_mem_slave_read -> NiosCustomIP2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nioscustomip2_debug_mem_slave_byteenable;  // mm_interconnect_0:NiosCustomIP2_debug_mem_slave_byteenable -> NiosCustomIP2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nioscustomip2_debug_mem_slave_write;       // mm_interconnect_0:NiosCustomIP2_debug_mem_slave_write -> NiosCustomIP2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nioscustomip2_debug_mem_slave_writedata;   // mm_interconnect_0:NiosCustomIP2_debug_mem_slave_writedata -> NiosCustomIP2:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                        // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                          // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [13:0] mm_interconnect_0_sram_s1_address;                           // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                        // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                             // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                         // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                             // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         irq_mapper_receiver0_irq;                                    // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nioscustomip2_irq_irq;                                       // irq_mapper:sender_irq -> NiosCustomIP2:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [DEBUG:rst_n, MyReg_0:reset_n, NiosCustomIP2:reset_n, SRAM:reset, irq_mapper:reset, mm_interconnect_0:NiosCustomIP2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [NiosCustomIP2:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	Nios_Custom_IP2_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	CustomIP myreg_0 (
		.address    (mm_interconnect_0_myreg_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_myreg_0_avalon_slave_0_chipselect), //               .chipselect
		.read       (mm_interconnect_0_myreg_0_avalon_slave_0_read),       //               .read
		.write      (mm_interconnect_0_myreg_0_avalon_slave_0_write),      //               .write
		.writedata  (mm_interconnect_0_myreg_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_myreg_0_avalon_slave_0_readdata),   //               .readdata
		.clk        (clk_clk),                                             //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset)                      //          reset.reset_n
	);

	Nios_Custom_IP2_NiosCustomIP2 nioscustomip2 (
		.clk                                 (clk_clk),                                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (nioscustomip2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nioscustomip2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nioscustomip2_data_master_read),                              //                          .read
		.d_readdata                          (nioscustomip2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nioscustomip2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nioscustomip2_data_master_write),                             //                          .write
		.d_writedata                         (nioscustomip2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nioscustomip2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nioscustomip2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nioscustomip2_instruction_master_read),                       //                          .read
		.i_readdata                          (nioscustomip2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nioscustomip2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nioscustomip2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nioscustomip2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nioscustomip2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nioscustomip2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nioscustomip2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nioscustomip2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nioscustomip2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nioscustomip2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nioscustomip2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nioscustomip2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                             // custom_instruction_master.readra
	);

	Nios_Custom_IP2_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	Nios_Custom_IP2_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                   (clk_clk),                                                     //                                 clk_0_clk.clk
		.NiosCustomIP2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // NiosCustomIP2_reset_reset_bridge_in_reset.reset
		.NiosCustomIP2_data_master_address               (nioscustomip2_data_master_address),                           //                 NiosCustomIP2_data_master.address
		.NiosCustomIP2_data_master_waitrequest           (nioscustomip2_data_master_waitrequest),                       //                                          .waitrequest
		.NiosCustomIP2_data_master_byteenable            (nioscustomip2_data_master_byteenable),                        //                                          .byteenable
		.NiosCustomIP2_data_master_read                  (nioscustomip2_data_master_read),                              //                                          .read
		.NiosCustomIP2_data_master_readdata              (nioscustomip2_data_master_readdata),                          //                                          .readdata
		.NiosCustomIP2_data_master_write                 (nioscustomip2_data_master_write),                             //                                          .write
		.NiosCustomIP2_data_master_writedata             (nioscustomip2_data_master_writedata),                         //                                          .writedata
		.NiosCustomIP2_data_master_debugaccess           (nioscustomip2_data_master_debugaccess),                       //                                          .debugaccess
		.NiosCustomIP2_instruction_master_address        (nioscustomip2_instruction_master_address),                    //          NiosCustomIP2_instruction_master.address
		.NiosCustomIP2_instruction_master_waitrequest    (nioscustomip2_instruction_master_waitrequest),                //                                          .waitrequest
		.NiosCustomIP2_instruction_master_read           (nioscustomip2_instruction_master_read),                       //                                          .read
		.NiosCustomIP2_instruction_master_readdata       (nioscustomip2_instruction_master_readdata),                   //                                          .readdata
		.DEBUG_avalon_jtag_slave_address                 (mm_interconnect_0_debug_avalon_jtag_slave_address),           //                   DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write                   (mm_interconnect_0_debug_avalon_jtag_slave_write),             //                                          .write
		.DEBUG_avalon_jtag_slave_read                    (mm_interconnect_0_debug_avalon_jtag_slave_read),              //                                          .read
		.DEBUG_avalon_jtag_slave_readdata                (mm_interconnect_0_debug_avalon_jtag_slave_readdata),          //                                          .readdata
		.DEBUG_avalon_jtag_slave_writedata               (mm_interconnect_0_debug_avalon_jtag_slave_writedata),         //                                          .writedata
		.DEBUG_avalon_jtag_slave_waitrequest             (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),       //                                          .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect              (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),        //                                          .chipselect
		.MyReg_0_avalon_slave_0_address                  (mm_interconnect_0_myreg_0_avalon_slave_0_address),            //                    MyReg_0_avalon_slave_0.address
		.MyReg_0_avalon_slave_0_write                    (mm_interconnect_0_myreg_0_avalon_slave_0_write),              //                                          .write
		.MyReg_0_avalon_slave_0_read                     (mm_interconnect_0_myreg_0_avalon_slave_0_read),               //                                          .read
		.MyReg_0_avalon_slave_0_readdata                 (mm_interconnect_0_myreg_0_avalon_slave_0_readdata),           //                                          .readdata
		.MyReg_0_avalon_slave_0_writedata                (mm_interconnect_0_myreg_0_avalon_slave_0_writedata),          //                                          .writedata
		.MyReg_0_avalon_slave_0_chipselect               (mm_interconnect_0_myreg_0_avalon_slave_0_chipselect),         //                                          .chipselect
		.NiosCustomIP2_debug_mem_slave_address           (mm_interconnect_0_nioscustomip2_debug_mem_slave_address),     //             NiosCustomIP2_debug_mem_slave.address
		.NiosCustomIP2_debug_mem_slave_write             (mm_interconnect_0_nioscustomip2_debug_mem_slave_write),       //                                          .write
		.NiosCustomIP2_debug_mem_slave_read              (mm_interconnect_0_nioscustomip2_debug_mem_slave_read),        //                                          .read
		.NiosCustomIP2_debug_mem_slave_readdata          (mm_interconnect_0_nioscustomip2_debug_mem_slave_readdata),    //                                          .readdata
		.NiosCustomIP2_debug_mem_slave_writedata         (mm_interconnect_0_nioscustomip2_debug_mem_slave_writedata),   //                                          .writedata
		.NiosCustomIP2_debug_mem_slave_byteenable        (mm_interconnect_0_nioscustomip2_debug_mem_slave_byteenable),  //                                          .byteenable
		.NiosCustomIP2_debug_mem_slave_waitrequest       (mm_interconnect_0_nioscustomip2_debug_mem_slave_waitrequest), //                                          .waitrequest
		.NiosCustomIP2_debug_mem_slave_debugaccess       (mm_interconnect_0_nioscustomip2_debug_mem_slave_debugaccess), //                                          .debugaccess
		.SRAM_s1_address                                 (mm_interconnect_0_sram_s1_address),                           //                                   SRAM_s1.address
		.SRAM_s1_write                                   (mm_interconnect_0_sram_s1_write),                             //                                          .write
		.SRAM_s1_readdata                                (mm_interconnect_0_sram_s1_readdata),                          //                                          .readdata
		.SRAM_s1_writedata                               (mm_interconnect_0_sram_s1_writedata),                         //                                          .writedata
		.SRAM_s1_byteenable                              (mm_interconnect_0_sram_s1_byteenable),                        //                                          .byteenable
		.SRAM_s1_chipselect                              (mm_interconnect_0_sram_s1_chipselect),                        //                                          .chipselect
		.SRAM_s1_clken                                   (mm_interconnect_0_sram_s1_clken)                              //                                          .clken
	);

	Nios_Custom_IP2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nioscustomip2_irq_irq)           //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nioscustomip2_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),          // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),      //          .reset_req
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_in1      (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

endmodule
