
module Nios_Buffer (
	clk_clk);	

	input		clk_clk;
endmodule
