// NiosInst.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module NiosInst (
		input  wire  clk_clk  // clk.clk
	);

	wire         nioscustominstr_debug_reset_request_reset;                                         // NiosCustomInstr:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] nioscustominstr_custom_instruction_master_result;                                  // NiosCustomInstr_custom_instruction_master_translator:ci_slave_result -> NiosCustomInstr:E_ci_combo_result
	wire         nioscustominstr_custom_instruction_master_readra;                                  // NiosCustomInstr:E_ci_combo_readra -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nioscustominstr_custom_instruction_master_a;                                       // NiosCustomInstr:E_ci_combo_a -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nioscustominstr_custom_instruction_master_b;                                       // NiosCustomInstr:E_ci_combo_b -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nioscustominstr_custom_instruction_master_c;                                       // NiosCustomInstr:E_ci_combo_c -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_c
	wire         nioscustominstr_custom_instruction_master_readrb;                                  // NiosCustomInstr:E_ci_combo_readrb -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_readrb
	wire         nioscustominstr_custom_instruction_master_estatus;                                 // NiosCustomInstr:E_ci_combo_estatus -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] nioscustominstr_custom_instruction_master_ipending;                                // NiosCustomInstr:E_ci_combo_ipending -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_ipending
	wire  [31:0] nioscustominstr_custom_instruction_master_datab;                                   // NiosCustomInstr:E_ci_combo_datab -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nioscustominstr_custom_instruction_master_dataa;                                   // NiosCustomInstr:E_ci_combo_dataa -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_dataa
	wire         nioscustominstr_custom_instruction_master_writerc;                                 // NiosCustomInstr:E_ci_combo_writerc -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_writerc
	wire   [7:0] nioscustominstr_custom_instruction_master_n;                                       // NiosCustomInstr:E_ci_combo_n -> NiosCustomInstr_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_result;        // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_result -> NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_result
	wire         nioscustominstr_custom_instruction_master_translator_comb_ci_master_readra;        // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_readra -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_a;             // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_a -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_b;             // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_b -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nioscustominstr_custom_instruction_master_translator_comb_ci_master_readrb;        // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_readrb -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_c;             // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_c -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nioscustominstr_custom_instruction_master_translator_comb_ci_master_estatus;       // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_estatus -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_ipending;      // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_ipending -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_datab;         // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_datab -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_dataa;         // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_dataa -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nioscustominstr_custom_instruction_master_translator_comb_ci_master_writerc;       // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_writerc -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nioscustominstr_custom_instruction_master_translator_comb_ci_master_n;             // NiosCustomInstr_custom_instruction_master_translator:comb_ci_master_n -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_result;         // NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_result -> NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_readra;         // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_readra -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_a;              // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_a -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_b;              // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_b -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_readrb -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_c;              // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_c -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_estatus -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_ipending -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_datab;          // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_datab -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_dataa -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_writerc -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_n;              // NiosCustomInstr_custom_instruction_master_comb_xconnect:ci_master0_n -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_result; // MyAnd:result -> NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_master_datab -> MyAnd:datab
	wire  [31:0] nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // NiosCustomInstr_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> MyAnd:dataa
	wire  [31:0] nioscustominstr_data_master_readdata;                                              // mm_interconnect_0:NiosCustomInstr_data_master_readdata -> NiosCustomInstr:d_readdata
	wire         nioscustominstr_data_master_waitrequest;                                           // mm_interconnect_0:NiosCustomInstr_data_master_waitrequest -> NiosCustomInstr:d_waitrequest
	wire         nioscustominstr_data_master_debugaccess;                                           // NiosCustomInstr:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosCustomInstr_data_master_debugaccess
	wire  [17:0] nioscustominstr_data_master_address;                                               // NiosCustomInstr:d_address -> mm_interconnect_0:NiosCustomInstr_data_master_address
	wire   [3:0] nioscustominstr_data_master_byteenable;                                            // NiosCustomInstr:d_byteenable -> mm_interconnect_0:NiosCustomInstr_data_master_byteenable
	wire         nioscustominstr_data_master_read;                                                  // NiosCustomInstr:d_read -> mm_interconnect_0:NiosCustomInstr_data_master_read
	wire         nioscustominstr_data_master_readdatavalid;                                         // mm_interconnect_0:NiosCustomInstr_data_master_readdatavalid -> NiosCustomInstr:d_readdatavalid
	wire         nioscustominstr_data_master_write;                                                 // NiosCustomInstr:d_write -> mm_interconnect_0:NiosCustomInstr_data_master_write
	wire  [31:0] nioscustominstr_data_master_writedata;                                             // NiosCustomInstr:d_writedata -> mm_interconnect_0:NiosCustomInstr_data_master_writedata
	wire  [31:0] nioscustominstr_instruction_master_readdata;                                       // mm_interconnect_0:NiosCustomInstr_instruction_master_readdata -> NiosCustomInstr:i_readdata
	wire         nioscustominstr_instruction_master_waitrequest;                                    // mm_interconnect_0:NiosCustomInstr_instruction_master_waitrequest -> NiosCustomInstr:i_waitrequest
	wire  [17:0] nioscustominstr_instruction_master_address;                                        // NiosCustomInstr:i_address -> mm_interconnect_0:NiosCustomInstr_instruction_master_address
	wire         nioscustominstr_instruction_master_read;                                           // NiosCustomInstr:i_read -> mm_interconnect_0:NiosCustomInstr_instruction_master_read
	wire         nioscustominstr_instruction_master_readdatavalid;                                  // mm_interconnect_0:NiosCustomInstr_instruction_master_readdatavalid -> NiosCustomInstr:i_readdatavalid
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;                              // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;                                // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest;                             // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;                                 // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;                                    // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;                                   // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;                               // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_nioscustominstr_debug_mem_slave_readdata;                        // NiosCustomInstr:debug_mem_slave_readdata -> mm_interconnect_0:NiosCustomInstr_debug_mem_slave_readdata
	wire         mm_interconnect_0_nioscustominstr_debug_mem_slave_waitrequest;                     // NiosCustomInstr:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosCustomInstr_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nioscustominstr_debug_mem_slave_debugaccess;                     // mm_interconnect_0:NiosCustomInstr_debug_mem_slave_debugaccess -> NiosCustomInstr:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nioscustominstr_debug_mem_slave_address;                         // mm_interconnect_0:NiosCustomInstr_debug_mem_slave_address -> NiosCustomInstr:debug_mem_slave_address
	wire         mm_interconnect_0_nioscustominstr_debug_mem_slave_read;                            // mm_interconnect_0:NiosCustomInstr_debug_mem_slave_read -> NiosCustomInstr:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nioscustominstr_debug_mem_slave_byteenable;                      // mm_interconnect_0:NiosCustomInstr_debug_mem_slave_byteenable -> NiosCustomInstr:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nioscustominstr_debug_mem_slave_write;                           // mm_interconnect_0:NiosCustomInstr_debug_mem_slave_write -> NiosCustomInstr:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nioscustominstr_debug_mem_slave_writedata;                       // mm_interconnect_0:NiosCustomInstr_debug_mem_slave_writedata -> NiosCustomInstr:debug_mem_slave_writedata
	wire         mm_interconnect_0_sram_s1_chipselect;                                              // mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	wire  [31:0] mm_interconnect_0_sram_s1_readdata;                                                // SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	wire  [13:0] mm_interconnect_0_sram_s1_address;                                                 // mm_interconnect_0:SRAM_s1_address -> SRAM:address
	wire   [3:0] mm_interconnect_0_sram_s1_byteenable;                                              // mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_s1_write;                                                   // mm_interconnect_0:SRAM_s1_write -> SRAM:write
	wire  [31:0] mm_interconnect_0_sram_s1_writedata;                                               // mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	wire         mm_interconnect_0_sram_s1_clken;                                                   // mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	wire         irq_mapper_receiver0_irq;                                                          // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nioscustominstr_irq_irq;                                                           // irq_mapper:sender_irq -> NiosCustomInstr:irq
	wire         rst_controller_reset_out_reset;                                                    // rst_controller:reset_out -> [DEBUG:rst_n, NiosCustomInstr:reset_n, SRAM:reset, irq_mapper:reset, mm_interconnect_0:NiosCustomInstr_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                                // rst_controller:reset_req -> [NiosCustomInstr:reset_req, SRAM:reset_req, rst_translator:reset_req_in]

	NiosInst_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	CustomInstr myand (
		.dataa  (nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // nios_custom_instruction_slave.dataa
		.datab  (nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //                              .datab
		.result (nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_result)  //                              .result
	);

	NiosInst_NiosCustomInstr nioscustominstr (
		.clk                                 (clk_clk),                                                       //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                               //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                            //                          .reset_req
		.d_address                           (nioscustominstr_data_master_address),                           //               data_master.address
		.d_byteenable                        (nioscustominstr_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nioscustominstr_data_master_read),                              //                          .read
		.d_readdata                          (nioscustominstr_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nioscustominstr_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nioscustominstr_data_master_write),                             //                          .write
		.d_writedata                         (nioscustominstr_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nioscustominstr_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nioscustominstr_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nioscustominstr_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nioscustominstr_instruction_master_read),                       //                          .read
		.i_readdata                          (nioscustominstr_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nioscustominstr_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nioscustominstr_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nioscustominstr_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nioscustominstr_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nioscustominstr_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nioscustominstr_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nioscustominstr_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nioscustominstr_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nioscustominstr_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nioscustominstr_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nioscustominstr_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nioscustominstr_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_combo_result                   (nioscustominstr_custom_instruction_master_result),              // custom_instruction_master.result
		.E_ci_combo_a                        (nioscustominstr_custom_instruction_master_a),                   //                          .a
		.E_ci_combo_b                        (nioscustominstr_custom_instruction_master_b),                   //                          .b
		.E_ci_combo_c                        (nioscustominstr_custom_instruction_master_c),                   //                          .c
		.E_ci_combo_dataa                    (nioscustominstr_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_combo_datab                    (nioscustominstr_custom_instruction_master_datab),               //                          .datab
		.E_ci_combo_estatus                  (nioscustominstr_custom_instruction_master_estatus),             //                          .estatus
		.E_ci_combo_ipending                 (nioscustominstr_custom_instruction_master_ipending),            //                          .ipending
		.E_ci_combo_n                        (nioscustominstr_custom_instruction_master_n),                   //                          .n
		.E_ci_combo_readra                   (nioscustominstr_custom_instruction_master_readra),              //                          .readra
		.E_ci_combo_readrb                   (nioscustominstr_custom_instruction_master_readrb),              //                          .readrb
		.E_ci_combo_writerc                  (nioscustominstr_custom_instruction_master_writerc)              //                          .writerc
	);

	NiosInst_SRAM sram (
		.clk        (clk_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_sram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_sram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_sram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_sram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_sram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_sram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_sram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze     (1'b0)                                  // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nioscustominstr_custom_instruction_master_translator (
		.ci_slave_dataa            (nioscustominstr_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nioscustominstr_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nioscustominstr_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nioscustominstr_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nioscustominstr_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nioscustominstr_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nioscustominstr_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nioscustominstr_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nioscustominstr_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nioscustominstr_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (nioscustominstr_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (nioscustominstr_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (nioscustominstr_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nioscustominstr_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nioscustominstr_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nioscustominstr_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nioscustominstr_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nioscustominstr_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nioscustominstr_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nioscustominstr_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_done       (),                                                                             //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                         //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                         //    (terminated)
		.ci_slave_multi_result     (),                                                                             //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                                  //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                     //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                     //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                                     //    (terminated)
		.multi_ci_master_clk       (),                                                                             //    (terminated)
		.multi_ci_master_reset     (),                                                                             //    (terminated)
		.multi_ci_master_clken     (),                                                                             //    (terminated)
		.multi_ci_master_reset_req (),                                                                             //    (terminated)
		.multi_ci_master_start     (),                                                                             //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                         //    (terminated)
		.multi_ci_master_dataa     (),                                                                             //    (terminated)
		.multi_ci_master_datab     (),                                                                             //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                         //    (terminated)
		.multi_ci_master_n         (),                                                                             //    (terminated)
		.multi_ci_master_readra    (),                                                                             //    (terminated)
		.multi_ci_master_readrb    (),                                                                             //    (terminated)
		.multi_ci_master_writerc   (),                                                                             //    (terminated)
		.multi_ci_master_a         (),                                                                             //    (terminated)
		.multi_ci_master_b         (),                                                                             //    (terminated)
		.multi_ci_master_c         ()                                                                              //    (terminated)
	);

	NiosInst_NiosCustomInstr_custom_instruction_master_comb_xconnect nioscustominstr_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nioscustominstr_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nioscustominstr_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nioscustominstr_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nioscustominstr_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nioscustominstr_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nioscustominstr_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nioscustominstr_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nioscustominstr_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nioscustominstr_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) nioscustominstr_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nioscustominstr_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nioscustominstr_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                                  // (terminated)
		.ci_master_readra    (),                                                                                  // (terminated)
		.ci_master_readrb    (),                                                                                  // (terminated)
		.ci_master_writerc   (),                                                                                  // (terminated)
		.ci_master_a         (),                                                                                  // (terminated)
		.ci_master_b         (),                                                                                  // (terminated)
		.ci_master_c         (),                                                                                  // (terminated)
		.ci_master_ipending  (),                                                                                  // (terminated)
		.ci_master_estatus   (),                                                                                  // (terminated)
		.ci_master_clk       (),                                                                                  // (terminated)
		.ci_master_clken     (),                                                                                  // (terminated)
		.ci_master_reset_req (),                                                                                  // (terminated)
		.ci_master_reset     (),                                                                                  // (terminated)
		.ci_master_start     (),                                                                                  // (terminated)
		.ci_master_done      (1'b0),                                                                              // (terminated)
		.ci_slave_clk        (1'b0),                                                                              // (terminated)
		.ci_slave_clken      (1'b0),                                                                              // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                              // (terminated)
		.ci_slave_reset      (1'b0),                                                                              // (terminated)
		.ci_slave_start      (1'b0),                                                                              // (terminated)
		.ci_slave_done       ()                                                                                   // (terminated)
	);

	NiosInst_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                     (clk_clk),                                                       //                                   clk_0_clk.clk
		.NiosCustomInstr_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                // NiosCustomInstr_reset_reset_bridge_in_reset.reset
		.NiosCustomInstr_data_master_address               (nioscustominstr_data_master_address),                           //                 NiosCustomInstr_data_master.address
		.NiosCustomInstr_data_master_waitrequest           (nioscustominstr_data_master_waitrequest),                       //                                            .waitrequest
		.NiosCustomInstr_data_master_byteenable            (nioscustominstr_data_master_byteenable),                        //                                            .byteenable
		.NiosCustomInstr_data_master_read                  (nioscustominstr_data_master_read),                              //                                            .read
		.NiosCustomInstr_data_master_readdata              (nioscustominstr_data_master_readdata),                          //                                            .readdata
		.NiosCustomInstr_data_master_readdatavalid         (nioscustominstr_data_master_readdatavalid),                     //                                            .readdatavalid
		.NiosCustomInstr_data_master_write                 (nioscustominstr_data_master_write),                             //                                            .write
		.NiosCustomInstr_data_master_writedata             (nioscustominstr_data_master_writedata),                         //                                            .writedata
		.NiosCustomInstr_data_master_debugaccess           (nioscustominstr_data_master_debugaccess),                       //                                            .debugaccess
		.NiosCustomInstr_instruction_master_address        (nioscustominstr_instruction_master_address),                    //          NiosCustomInstr_instruction_master.address
		.NiosCustomInstr_instruction_master_waitrequest    (nioscustominstr_instruction_master_waitrequest),                //                                            .waitrequest
		.NiosCustomInstr_instruction_master_read           (nioscustominstr_instruction_master_read),                       //                                            .read
		.NiosCustomInstr_instruction_master_readdata       (nioscustominstr_instruction_master_readdata),                   //                                            .readdata
		.NiosCustomInstr_instruction_master_readdatavalid  (nioscustominstr_instruction_master_readdatavalid),              //                                            .readdatavalid
		.DEBUG_avalon_jtag_slave_address                   (mm_interconnect_0_debug_avalon_jtag_slave_address),             //                     DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write                     (mm_interconnect_0_debug_avalon_jtag_slave_write),               //                                            .write
		.DEBUG_avalon_jtag_slave_read                      (mm_interconnect_0_debug_avalon_jtag_slave_read),                //                                            .read
		.DEBUG_avalon_jtag_slave_readdata                  (mm_interconnect_0_debug_avalon_jtag_slave_readdata),            //                                            .readdata
		.DEBUG_avalon_jtag_slave_writedata                 (mm_interconnect_0_debug_avalon_jtag_slave_writedata),           //                                            .writedata
		.DEBUG_avalon_jtag_slave_waitrequest               (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest),         //                                            .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect                (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),          //                                            .chipselect
		.NiosCustomInstr_debug_mem_slave_address           (mm_interconnect_0_nioscustominstr_debug_mem_slave_address),     //             NiosCustomInstr_debug_mem_slave.address
		.NiosCustomInstr_debug_mem_slave_write             (mm_interconnect_0_nioscustominstr_debug_mem_slave_write),       //                                            .write
		.NiosCustomInstr_debug_mem_slave_read              (mm_interconnect_0_nioscustominstr_debug_mem_slave_read),        //                                            .read
		.NiosCustomInstr_debug_mem_slave_readdata          (mm_interconnect_0_nioscustominstr_debug_mem_slave_readdata),    //                                            .readdata
		.NiosCustomInstr_debug_mem_slave_writedata         (mm_interconnect_0_nioscustominstr_debug_mem_slave_writedata),   //                                            .writedata
		.NiosCustomInstr_debug_mem_slave_byteenable        (mm_interconnect_0_nioscustominstr_debug_mem_slave_byteenable),  //                                            .byteenable
		.NiosCustomInstr_debug_mem_slave_waitrequest       (mm_interconnect_0_nioscustominstr_debug_mem_slave_waitrequest), //                                            .waitrequest
		.NiosCustomInstr_debug_mem_slave_debugaccess       (mm_interconnect_0_nioscustominstr_debug_mem_slave_debugaccess), //                                            .debugaccess
		.SRAM_s1_address                                   (mm_interconnect_0_sram_s1_address),                             //                                     SRAM_s1.address
		.SRAM_s1_write                                     (mm_interconnect_0_sram_s1_write),                               //                                            .write
		.SRAM_s1_readdata                                  (mm_interconnect_0_sram_s1_readdata),                            //                                            .readdata
		.SRAM_s1_writedata                                 (mm_interconnect_0_sram_s1_writedata),                           //                                            .writedata
		.SRAM_s1_byteenable                                (mm_interconnect_0_sram_s1_byteenable),                          //                                            .byteenable
		.SRAM_s1_chipselect                                (mm_interconnect_0_sram_s1_chipselect),                          //                                            .chipselect
		.SRAM_s1_clken                                     (mm_interconnect_0_sram_s1_clken)                                //                                            .clken
	);

	NiosInst_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nioscustominstr_irq_irq)         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nioscustominstr_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),            // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),        //          .reset_req
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_in1      (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

endmodule
