
module nios_custom_dma (
	clk_clk);	

	input		clk_clk;
endmodule
