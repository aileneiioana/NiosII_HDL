	component acc_spi is
		port (
			accelerometer_spi_0_external_interface_I2C_SDAT      : inout std_logic := 'X'; -- I2C_SDAT
			accelerometer_spi_0_external_interface_I2C_SCLK      : out   std_logic;        -- I2C_SCLK
			accelerometer_spi_0_external_interface_G_SENSOR_CS_N : out   std_logic;        -- G_SENSOR_CS_N
			accelerometer_spi_0_external_interface_G_SENSOR_INT  : in    std_logic := 'X'; -- G_SENSOR_INT
			clk_clk                                              : in    std_logic := 'X'  -- clk
		);
	end component acc_spi;

	u0 : component acc_spi
		port map (
			accelerometer_spi_0_external_interface_I2C_SDAT      => CONNECTED_TO_accelerometer_spi_0_external_interface_I2C_SDAT,      -- accelerometer_spi_0_external_interface.I2C_SDAT
			accelerometer_spi_0_external_interface_I2C_SCLK      => CONNECTED_TO_accelerometer_spi_0_external_interface_I2C_SCLK,      --                                       .I2C_SCLK
			accelerometer_spi_0_external_interface_G_SENSOR_CS_N => CONNECTED_TO_accelerometer_spi_0_external_interface_G_SENSOR_CS_N, --                                       .G_SENSOR_CS_N
			accelerometer_spi_0_external_interface_G_SENSOR_INT  => CONNECTED_TO_accelerometer_spi_0_external_interface_G_SENSOR_INT,  --                                       .G_SENSOR_INT
			clk_clk                                              => CONNECTED_TO_clk_clk                                               --                                    clk.clk
		);

