
module Nios_Custom_IP2 (
	clk_clk);	

	input		clk_clk;
endmodule
