
module dma (
	clk_clk);	

	input		clk_clk;
endmodule
